-- --------------------------------------------------------------------
-- comp_pack.vhd
-- --------------------------------------------------------------------
-- FPGA-chip: 10M16SAU169C8G (most likely)  
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- last edited: 2020-0617
-- --------------------------------------------------------------------

LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.all;
  USE IEEE.NUMERIC_STD.all;

-- --------------------------------------------------------------------

PACKAGE comp_pack IS

COMPONENT top IS
PORT();
END COMPONENT;

END comp_pack;