ARCHITECTURE top_a OF top_e is
BEGIN



END top_a;