ARCHITECTURE rtc_a OF rtc_e is
BEGIN



END rtc_a;