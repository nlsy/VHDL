ARCHITECTURE uat_a OF uat_e is
BEGIN



END uat_a;